`include "define.v"

module fetch(clk, pc, instr);
	input clk;
	input pc;