`include "define.v"

module RRS();
endmodule